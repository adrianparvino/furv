(*blackbox*)
module rom(
  input [31:0] pc,
  output [31:0] instruction
);

endmodule
